----------------------------------------------------------------------------------------------------
--											inverter_maia_2.vhd										 ---
----------------------------------------------------------------------------------------------------
--	Inverter for F_2^m 
----------------------------------------------------------------------------------------------------
-- Author		: Miguel Morales-Sandoval														 ---
-- Project		: "Hardware Arquitecture for ECC and Lossless Data Compression					 ---
-- Organization	: INAOE, Computer Science Department											 ---
-- Date			: July, 2004.																	 ---
----------------------------------------------------------------------------------------------------
-- Coments: This is an implementation of the Modified Almost Inverse Algorithm.
--			Diferent to the first implementation, here the test g(U) < g(V) is
--			performed directly by a m+1 bit comparer.
----------------------------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all; 
use IEEE.STD_LOGIC_unsigned.all; 
use IEEE.STD_LOGIC_arith.all;
--------------------------------------------------------
entity inverter_maia_163 is
	generic(       
		NUM_BITS : positive := 163							-- The order of the finite field
	);
	port( 
		 ax    : in STD_LOGIC_VECTOR(NUM_BITS-1 downto 0); 	-- input polynomial of grade m-1
		 clk  : in STD_LOGIC;
		 rst  : in STD_LOGIC;
		 done : out STD_LOGIC;
		 z    : out STD_LOGIC_VECTOR(NUM_BITS-1 downto 0)
	     );
end ;
---------------------------------------------------------
architecture behave of inverter_maia_163 is		
---------------------------------------------------------
	signal B,C,U,V  : STD_LOGIC_VECTOR(NUM_BITS downto 0);  -- Internal processing registers, one bit more
	signal Bx_Op1   : STD_LOGIC_VECTOR(NUM_BITS downto 0);  -- Multiplexer which depends on if B is ever or odd
	signal Ux_div_x : STD_LOGIC_VECTOR(NUM_BITS downto 0);  -- U and B divided by x
	signal Bx_div_x : STD_LOGIC_VECTOR(NUM_BITS downto 0);  
	--163
	constant UNO    : STD_LOGIC_VECTOR(NUM_BITS downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";															  
	--233
--	constant UNO    : STD_LOGIC_VECTOR(NUM_BITS downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";
	--277
--	constant UNO    : STD_LOGIC_VECTOR(NUM_BITS downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";
	--283
--	constant UNO    : STD_LOGIC_VECTOR(NUM_BITS downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";
	--409
--	constant UNO    : STD_LOGIC_VECTOR(NUM_BITS downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";
	--571
--	constant UNO    : STD_LOGIC_VECTOR(NUM_BITS downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";
--	
-- m = 163		  x163 + x7 + x6 + x3 + 1
constant Fx: std_logic_vector(NUM_BITS downto 0) := "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001";
-- m = 233		  x233 + x74 + 1
--constant Fx: std_logic_vector(NUM_BITS downto 0) := "100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000001";
-- m = 277		  x277 + x74 + 1
--constant Fx: std_logic_vector(NUM_BITS downto 0) := "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001001001"; --277 bits
-- m = 283        x283 + x12 + x7 + x5 + 1														
--constant Fx: std_logic_vector(NUM_BITS downto 0) := "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010100001";
-- m = 409		  x409 + x87 + 1
--constant Fx: std_logic_vector(NUM_BITS1 downto 0) := "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";
-- m = 571        x571 + x10 + x5 + x2 + 1													
--constant Fx: std_logic_vector(NUM_BITS downto 0) := "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100101";

	----------------------------------------------------------------------------------
	-- States fot the FSM controlling the execution of the algorithm
	----------------------------------------------------------------------------------
	type CurrentState_type is (END_STATE, LOOP_U0, NEXT_STEP);
	signal State: CurrentState_type;
	----------------------------------------------------------------------------------
begin			  
	
	------------------------------------------------------
	Ux_div_x <= '0' & U(NUM_BITS downto 1);					-- Dividing U and B by x
	Bx_div_x <= '0' & Bx_Op1(NUM_BITS downto 1);
	------------------------------------------------------
	Bx_Op1   <= B xor Fx when B(0) = '1' else				-- Multiplexer for operand B 
		        B;
	-------------------------------------------------------
	-- The Modified ALmost Inverse Algorithm implementation
	-------------------------------------------------------
	EEAL: process (clk)
		begin -- syncronous reset
			if CLK'event and CLK = '1' then
				if (rst = '1')then							-- initialize internal registers
					State <= LOOP_U0;	 	
					B <= UNO;
					U <= '0'&Ax;
					V <= Fx;
					C <= (others => '0');					
					z <= (others => '0');					-- set to zero the output register
					Done      <= '0';					
				else	
					case State is 
						-----------------------------------------------------------------------------------
						when LOOP_U0 =>						-- Stay here while U be even
							if U(0) = '1' then
								if U = UNO then				-- The algorithm finishes when U = 1
									Z <= B(NUM_BITS-1 downto 0);
									Done <= '1';
									State <= END_STATE;
								else						
									if U < V then			-- Interchange the registers U <-> V and B <-> C
										U <= V;
										V <= U;
										B <= C;
										C <= B;
									end if;	   
									
									State <= NEXT_STEP;	
								end if;
							else							-- Divide U and B and repeat the process
								U <= Ux_div_x;
								B <= Bx_div_x;
							end if;
						-----------------------------------------------------------------------------------	
						when NEXT_STEP => 					-- update U and B with the values previously assigned
							U <= U xor V;
							B <= B xor C;
							State <= LOOP_U0;
						 -----------------------------------------------------------------------------------
						when END_STATE =>					-- Do nothing 
							State <= END_STATE;
						-----------------------------------------------------------------------------------
						when others =>
							null;
					end case;
				end if;
			end if;			
		end process;
end behave;